`define DIV
