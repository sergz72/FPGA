`define STAGE_WIDTH 2
//`define NO_MUL
//`define NO_DIV
