//`define NO_MUL
`define NO_DIV1616
`define NO_REM1616
`define NO_DIV3216
`define NO_REM3216
