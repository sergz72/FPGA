`define ALU_OP_TEST  0
`define ALU_OP_NOT   1
`define ALU_OP_NEG   2
`define ALU_OP_ADD   3
`define ALU_OP_ADC   4
`define ALU_OP_SUB   5
`define ALU_OP_SBC   6
`define ALU_OP_SHL   7
`define ALU_OP_SHR   8

`define ALU_OPID_WIDTH 5
