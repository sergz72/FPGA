//`define NO_MUL
`define NO_DIV
`define NO_REM
