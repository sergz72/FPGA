//`define INTEL
