`define ALU_OP_NOP   0
`define ALU_OP_ZERO  1
`define ALU_OP_NZERO 2
`define ALU_OP_TEST  3
`define ALU_OP_NOT   4
`define ALU_OP_NEG   5
`define ALU_OP_INC   6
`define ALU_OP_DEC   7
`define ALU_OP_ADD   8
`define ALU_OP_ADC   9
`define ALU_OP_SUB   10
`define ALU_OP_SBC   11
`define ALU_OP_SHL   12
`define ALU_OP_SHR   13

`define ALU_OPID_WIDTH 5
