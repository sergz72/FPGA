`define STAGE_WIDTH 3
//`define NO_MUL
//`define NO_DIV
