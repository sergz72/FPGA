`define DIV
`define REM
