//`define MUL
