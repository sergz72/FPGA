`define MEMORY_DEBUG
