`define ALU_OP_TEST  0
`define ALU_OP_CMP   1
`define ALU_OP_SETF  2

`define ALU_OP_NEG   4
`define ALU_OP_ADD   5
`define ALU_OP_ADC   6
`define ALU_OP_SUB   7
`define ALU_OP_SBC   8
`define ALU_OP_SHL   9
`define ALU_OP_SHR   10
`define ALU_OP_AND   11
`define ALU_OP_OR    12
`define ALU_OP_XOR   13
`define ALU_OP_RLC   14
`define ALU_OP_RRC   15
`define ALU_OP_SHLC  16
`define ALU_OP_SHRC  17

`define ALU_OP_DIV1616   27
`define ALU_OP_REM1616   28
`define ALU_OP_DIV3216   29
`define ALU_OP_REM3216   30
`define ALU_OP_MUL       31

`define ALU_OPID_WIDTH 5
