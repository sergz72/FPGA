`define STAGE_WIDTH 3
`define DIV
`define REM
