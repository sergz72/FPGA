`define MEMORY_DEBUG
