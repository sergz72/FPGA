`define NO_DIV
`define NO_REM
`define NO_MUL
