`define MEMORY_DEBUG
`define UART_CLOCK_DIV 8
`define UART_CLOCK_COUNTER_BITS 4
`define CPU_TIMER_BITS 6
`define CPU_CLOCK_BIT 3
`define MHZ_TIMER_BITS 1
`define MHZ_TIMER_VALUE 1
