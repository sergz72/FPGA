`define NO_DIV
`define NO_REM
