`define CPU_TIMER_BITS 3
`define CPU_CLOCK_BIT 0
`define MHZ_TIMER_BITS 1
`define MHZ_TIMER_VALUE 1
