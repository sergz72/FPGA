//`define MUL
//`define loadpc
