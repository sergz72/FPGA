`define RAM
`define CHARACTER_ROM
