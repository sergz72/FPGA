//`define DIV
