//`define RAM
//`define CHARACTER_ROM
`define INTEL
