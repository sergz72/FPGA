`define MEMORY_DEBUG
`define OSC_FREQ 2000000
