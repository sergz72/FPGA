//`define NO_MUL
//`define NO_DIV
