//`define MUL
//`define DIV
