`define MUL
`define DIV
