`define QSPI_DATA_8_15
`define QSPI_DATA_16_31
