`define ALU_OP_TEST  0
`define ALU_OP_NEG   1
`define ALU_OP_ADD   2
`define ALU_OP_ADC   3
`define ALU_OP_SUB   4
`define ALU_OP_SBC   5
`define ALU_OP_SHL   6
`define ALU_OP_SHR   7
`define ALU_OP_AND   8
`define ALU_OP_OR    9
`define ALU_OP_XOR   10
`define ALU_OP_CMP   11
`define ALU_OP_MUL   12
`define ALU_OP_DIV   13
`define ALU_OP_REM   14
`define ALU_OP_SETF  15

`define ALU_OPID_WIDTH 5
