`define CPU_TIMER_BITS 3
`define CPU_CLOCK_BIT 0
