`define NO_DIV
`define NO_MUL
