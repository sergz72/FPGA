//`define NO_DIV
